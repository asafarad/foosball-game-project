//-- Alex Grinshpun Apr 2017
//-- Dudy Nov 13 2017
// SystemVerilog version Alex Grinshpun May 2018



module	ball_object	(	
//		--////////////////////	Clock Input	 	////////////////////	
					input		logic	CLK,
					input		logic	RESETn,
					input 	logic	[10:0]	oCoord_X,
					input 	logic	[10:0]	oCoord_Y,
					input 	logic	[10:0]	ObjectStartX,
					input 	logic	[10:0]	ObjectStartY,
					input		logic 			double_ball_ena,
					output	logic				drawing_request,
					output	logic	[7:0]		mVGA_RGB
					
);

localparam  int object_X_size = 26;
localparam  int object_Y_size = 26;


bit [0:object_Y_size-1] [0:object_X_size-1] [7:0] object_colors = {
{8'h00,8'h00,8'h00,8'h92,8'h92,8'h6d,8'hb6,8'h49,8'h00,8'h00,8'h49,8'h49,8'h92,8'hb6,8'hb6,8'h6d,8'h00,8'h00,8'h6d,8'hdb,8'h6d,8'h92,8'h92,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h49,8'h49,8'h49,8'h92,8'hdb,8'hdb,8'hdb,8'hdb,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h92,8'h49,8'h49,8'hb6,8'hb6,8'hdb,8'hdb,8'h00,8'h00},
{8'h00,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hb6,8'h92,8'h24,8'h6d,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hb6,8'h00,8'h00,8'h92,8'hdb,8'hb6,8'h00},
{8'h92,8'h92,8'h6d,8'h49,8'h49,8'h49,8'h24,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h49,8'h49,8'h92,8'h92,8'h92},
{8'h49,8'h92,8'hff,8'hdb,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h49,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h92,8'h00,8'hb6,8'hff,8'h49,8'h49,8'h92,8'h49},
{8'h6d,8'h6d,8'h49,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h24,8'h00,8'h00,8'h00,8'hb6,8'hff,8'h00,8'h00,8'h6d},
{8'hff,8'hff,8'hdb,8'h92,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hdb,8'hff,8'hff},
{8'h6d,8'h49,8'hff,8'h6d,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hdb,8'h6d,8'h92},
{8'hff,8'hdb,8'hff,8'hdb,8'hb6,8'hb6,8'h92,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hff},
{8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'h00},
{8'h92,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h49,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'h6d},
{8'h92,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hff,8'hff,8'hb6,8'h6d,8'h92,8'hff,8'hff,8'h92},
{8'h49,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6},
{8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6},
{8'h00,8'h92,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h6d,8'h00,8'h24,8'h49,8'h6d,8'hb6,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h92},
{8'h00,8'h49,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h6d},
{8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hdb,8'h00},
{8'h00,8'h00,8'h6d,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h24,8'h24},
{8'h00,8'h00,8'h6d,8'hff,8'hdb,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h24,8'h00,8'h00,8'h00},
{8'hff,8'hff,8'h6d,8'hff,8'hff,8'hff,8'hff,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'h49,8'h00,8'h00,8'h00,8'h00},
{8'h92,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00,8'h92,8'hff,8'hdb,8'hff,8'hff,8'hdb,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h92,8'h92,8'h6d,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h6d,8'h00,8'h49,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h92,8'h92,8'h92,8'h49,8'h6d,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'hb6,8'hdb,8'h92,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'hdb,8'hdb,8'hb6,8'hdb,8'hdb,8'h6d,8'hb6,8'h92,8'h92,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h6d,8'h92,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00},
{8'h00,8'h00,8'h00,8'h92,8'h92,8'h6d,8'hdb,8'h49,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hb6,8'hb6,8'h6d,8'h00,8'h00,8'hdb,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}
};

//-- one bit mask  0 - off 1 dispaly 

bit [0:object_Y_size-1] [0:object_X_size-1] object_mask = {
{26'b00000000000000000000000000},
{26'b00000011111111111111000000},
{26'b00000111111111111111100000},
{26'b00001111111111111111110000},
{26'b00011111111111111111111000},
{26'b00111111111111111111111100},
{26'b00111111111111111111111110},
{26'b01111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b11111111111111111111111111},
{26'b01111111111111111111111110},
{26'b00111111111111111111111100},
{26'b00011111111111111111111000},
{26'b00001111111111111111110000},
{26'b00000111111111111111100000},
{26'b00000011111111111111000000},
{26'b00000000000000000000000000}
};   
  

int bCoord_X ;// offset from start position 
int bCoord_Y ;

logic drawing_X ;  /* synthesis keep */
logic drawing_Y ; /* synthesis keep */
logic mask_bit	; /* synthesis keep */

int objectEndX ;
int objectEndY ;



// Calculate object end boundaries
assign objectEndX	= (object_X_size + ObjectStartX);
assign objectEndY	= (object_Y_size + ObjectStartY);
//
//-- Signals drawing_X[Y] are active when obects coordinates are being crossed
//
//-- test if ooCoord is in the rectangle defined by Start and End 

assign drawing_X	= ((oCoord_X  >= ObjectStartX) &&  (oCoord_X < objectEndX)) ? 1 : 0;
assign drawing_Y	= ((oCoord_Y  >= ObjectStartY) &&  (oCoord_Y < objectEndY)) ? 1 : 0;

assign bCoord_X	= (drawing_X == 1 &&  drawing_Y == 1  )  ? (oCoord_X - ObjectStartX): 0;
assign bCoord_Y	= (drawing_X == 1 &&  drawing_Y == 1  )  ? (oCoord_Y - ObjectStartY): 0;



always_ff@(posedge CLK or negedge RESETn)
begin
	if(!RESETn)
	begin
		mVGA_RGB				<=	8'b0;
		drawing_request	<=	1'b0;
		mask_bit				<=	1'b0;
	end
	else
	begin
		mVGA_RGB				<= object_colors[bCoord_Y][bCoord_X];	//get from colors table 
		drawing_request	<= object_mask[bCoord_Y][bCoord_X] && drawing_X && drawing_Y && double_ball_ena; // get from mask table if inside rectangle and enable
		mask_bit				<= object_mask[bCoord_Y][bCoord_X];
	end
end



endmodule