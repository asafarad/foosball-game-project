module game_over_object (
	   	input   logic   CLK,
		input   logic   RESETn,
		input   logic [10:0] oCoord_X,
		input   logic [10:0] oCoord_Y,
		input   logic game_over_ena,
		output  logic   drawing_request,		
		output  logic [7:0] mVGA_RGB 
);

localparam int object_X_size = 120;
localparam int object_Y_size = 120;


// one bit mask  0 - off 1 dispaly 
bit [0:object_Y_size-1] [0:object_X_size-1] object_mask = {
{120'b000000000001100000000000110000000000000000000000000000000001011111110100000000000001011100000000000000000000000000000000},
{120'b000000000010111111111111101000000000000000000000000000000001011111110100000000000010111100000000000000000000000000000000},
{120'b000000000010111111111111110100000000000000000000000000000001011111111010000000000010111100000000000000000000000000000000},
{120'b000000000101111111111111111010000000000000000000000000000001011111111010000000000101111100000000000000000000000000000010},
{120'b000000001011111111111111111101000000000000000110000000000001011111111101000000000101111100000000000000000000000000111100},
{120'b000000001011111111111111111110100000000000001010000000000001011111111101000000001011111100000000000000000000000111000010},
{120'b000000010111111111111111111110100000000000010110000000000001011111111110100000001011111100000000000000000001111000111111},
{120'b000000010111111111111111111110100000000000101110100000000001011111111110100000010111111101000000000000001110000111111111},
{120'b000000101111111111111111111110100000000000011111010000000001011111111110100000010111111101000000000011110001111111111111},
{120'b000000101111111111111111111110100000000001011111101000000001011111111111010000101111111101000000011100001111111111111111},
{120'b000001011111111111111111111110100000000010111111101000000001011111111111010000101111111101000111000011111111111111111111},
{120'b000001011111111111111111111110100000000010111111110100000001011111111111101001011111111101011001011111111111111111111111},
{120'b000010111111111111111111111110100000000101111111110100000001011111111111101001011111111101100111111111111111111111111111},
{120'b000010111111111111111111111110100000000101111111111010000001011111111111110110111111111101111111111111111111111111111111},
{120'b000101111111111110111111111110100000001011111111111101000001011111111111110110111111111101111111111111111111111111111111},
{120'b001011111111111110101111111110100000010111111111111101000001011111111111111001111111111101111111111111111111111111111111},
{120'b001011111111111101110111111110100000010111111111111110100001011111111111111111111111111101111111111111111111111111111111},
{120'b010111111111111101011101111110100000101111111111111111010001011111111111111111111111111101111111111111111111111111111111},
{120'b010111111111111010000110001110000000101111111111111111010001011111111111111111111111111101111111111111111111111111111111},
{120'b101111111111111010000001110000000001011111111111111111101001011111111111111111111111111101111111111111111111111111111111},
{120'b101111111111110100000000001100000001011111111111111111101001011111111111111111111111111101111111111111111111111111111111},
{120'b011111111111110100000000000111000010111111111111111111110101011111111111111111111111111101111111111111111111111111111111},
{120'b011111111111101001111111100000000010111111111111111111111011011111111111111111111111111101111111111111111111111111111111},
{120'b111111111111101000000000011111100101111111111111111111111011011111111111111111111111111101111111111111111111111111111111},
{120'b111111111111010101111111111111101101111111111111111111111101011111111111111111111111111101111111111111111111111111111110},
{120'b111111111111010101111111111111101101111111111111111111111110011111111111111111111111111101111111111111111111111111110000},
{120'b111111111111010101111111111111101101111111111111111111111110011111111111111111111111111101111111111111111111111000000000},
{120'b111111111111010101111111111111101011111111111111111111111110011111111111111111111111111101111111111111111100000000000000},
{120'b111111111111010101111111111111101011111111111111111111111110011111111111111111111111111101111111111111111111110000000000},
{120'b111111111111010101111111111111101011111111111111111111111110011111111111111111111111111101111111111111111111111110000000},
{120'b111111111111010101111111111111101011111111111111111111111110011111111111111111111111111101111111111111111111111111000000},
{120'b111111111111010101111111111111101011111111111101111111111110011111111111111111111111111101111111111111111111111111000000},
{120'b111111111111010101111111111111100111111111110001111111111110011111111111111111111111111101111111111111111111111111000000},
{120'b111111111111010101111111111111100111111111110000111111111111001111111111111111111111111101111111111111111111111111000000},
{120'b111111111111010000001111111111100111111111110001111111111110011111111111111111111111111101111111111111111111111111000000},
{120'b111111111111010001110101111111100111111111110001111111111110011111111111111111111111111101111111111111111111111111000000},
{120'b111111111111101100011101111111101111111111110001111111111110011111111111111111111111111101111111111111111111111111000000},
{120'b111111111111110111111101111111101111111111110001111111111110011111111111111111111111111101111111111111111111111111000000},
{120'b111111111111111101000101111111101111111111111111111111111110011111111111111111111111111101111111111111111111111111000000},
{120'b111111111111111111111111111111101111111111111111111111111110011111111111111111110111111101111111111111111111111110000000},
{120'b111111111111111111111111111111101111111111111111111111111110011111111111111111110111111101111111111111111111111110000000},
{120'b111111111111111111111111111111111111111111111111111111111110111111111111111111110111111101111111111111111111110000000000},
{120'b111111111111111111111111111111111111111111111111111111111110111111111101111111100111111101111111111111111110100000000000},
{120'b111111111111111111111111111111111111111111111111111111111110111111111101111111010111111101111111111111110000000000000000},
{120'b111111111111111111111111111111111111111111111111111111111110111111111101111111010111111101111111111111110000000000000000},
{120'b111111111111111111111111111111111111111111111111111111111110111111111100111110110111111101111111111111111111111111111000},
{120'b011111111111111111111111111111111111111111111111111111111110111111111100111110110111111101111111111111111111111111111101},
{120'b011111111111111111111111111111111111111111111111111111111110111111111100111101010111111101111111111111111111111111111101},
{120'b101111111111111111111111111111111111111111111111111111111110111111111001011101010111111101111111111111111111111111111101},
{120'b101111111111111111111111111111111111111111111111111111111111111111111011011101010111111101111111111111111111111111111101},
{120'b010111111111111111111111111111111111111111111111111111111111111111111010011000010111111101111111111111111111111111111101},
{120'b001011111111111111111111111111111111111111111111111111111111111111111010001100010111111101111111111111111111111111111101},
{120'b001011111111111111111111111101111111111111111011111111111111111111111010001000010111111101111111111111111111111111111101},
{120'b000101111111111111111111111101111111111111101011111111111111111111111010000000010111111101111111111111111111111111111101},
{120'b000101111111111111111111111111111111111111101011111111111111111111111010000000010111111101111111111111111111111111111101},
{120'b000010111111111111111111111011111111111111011011111111111111111111111010000000010111111101111111111111111111111111111101},
{120'b000010111111111111111111111011111111111111011011111111111111111111111010000000010111111101111111111111111111111111111101},
{120'b000001011111111111111111111011111111111111011011111111111111111111110000000000010111111101101111111111111111111111111101},
{120'b000000101111111111111111110011111111111110101011111111111111111111110100000000000111111101101111111111111111111111111101},
{120'b000000101111111111111111110100000000000100000001111111111110011111110000000000000100000000001111111111111111111111111100},
{120'b000000001010111111111010010011111110111110100010000000000001100000000000000001111000111110100000000000000000011101000000},
{120'b000000001101111111111011110000111011111110100101110111111100011111100000000110010111111110101111111111111001111101111000},
{120'b000000000101111111111101000001101111111110100101111010000000000000000011110001111111111110100000000111101111111110100000},
{120'b000000001011111111111110100010111111111110010101111101000000000000011110001111111111111110100000001100111111111110100000},
{120'b000000001011111111111110100101111111111111010101111110100000000111100011111111111111111110100001100111111111111111010000},
{120'b000000010111111111111111011011111111111111010101111111010000111100011111111111111111111110100111011111111111111111101000},
{120'b000000010111111111111111011011111111111111010101111111101011000111111111111111111111111110111101111111111111111111101000},
{120'b000000101111111111111111101011111111111111010101111111110100111111111111111111111111111110110111111111111111111111110100},
{120'b000001011111111111111111101101111111111111010101111111111011111111111111111111111111111110011111111111111111111111110100},
{120'b000001011111111111111111110101111111111111011011111111111011111111111111111111111111111110111111111111111111111111111010},
{120'b000010111111111111111111111001111111111111101011111111111111111111111111111111111111111111111111111111111111111111111010},
{120'b000010111111111111111111111001111111111111101011111111111111111111111111111111111111111111111111111111111111111111111101},
{120'b000101111111111111111111111100111111111111101011111111111111111111111111111111111111111111111111111111111111111111111101},
{120'b000101111111111111111111111100111111111111101011111111111111111111111111111111111111111111111111111111111111111111111110},
{120'b001011111111111111111111111110111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111},
{120'b001011111111111101111111111111111111111111101011111111111111111111111111111111111111111111111111111111111111111111111111},
{120'b010111111111111100111111111111011111111111101011111111111111111111111111111111111111111111111111111111111111111111111111},
{120'b010111111111111010111111111111111111111111101011111111111101111111111111111111111111111111111111111111111111111111111111},
{120'b101111111111111010111111111111111111111111110011111111111101111111111111111111111111111111111111111111011111111111111111},
{120'b101111111111110110011111111111111111111111110011111111111101111111111111111111111111111101111111111111001111111111111111},
{120'b011111111111110101011111111111101111111111110011111111111101111111111111111111111100000101111111111111010111111111111111},
{120'b011111111111101001011111111111101111111111110011111111111101111111111111111110000111111101111111111111011011111111111111},
{120'b111111111111100001011111111111101111111111110111111111111001111111111111111101000000000101111111111111010101111111111111},
{120'b111111111111010000101111111111101111111111110111111111111001111111111111111111111110100101111111111111010101111111111111},
{120'b111111111111010000101111111111101111111111110111111111111001111111111111111111111110100101111111111111010101111111111111},
{120'b111111111111010000101111111111100111111111110111111111111001111111111111111111111110100101111111111111010101111111111111},
{120'b111111111111101001011111111111100111111111111111111111110101111111111111111111111110100101111111111111010101111111111111},
{120'b111111111111101001011111111111100111111111111111111111110101111111111111111111111110100101111111111111010101111111111111},
{120'b111111111111110101011111111111100111111111111111111111110101111111111111111111111110100101111111111111010101111111111110},
{120'b111111111111110110111111111111101011111111111111111111110101111111111111111111111110100101111111111111010101111111111110},
{120'b111111111111111010111111111111101011111111111111111111110101111111111111111111111110100101111111111111010101111111111101},
{120'b111111111111111110111111111111101011111111111111111111101101111111111111111111111110100101111111111111011101111111111010},
{120'b111111111111111101111111111111101011111111111111111111101100111111111111111111111110100101111111111111011011111111111010},
{120'b111111111111111111111111111111101101111111111111111111101010111111111111111111111110100101111111111111011111111111110100},
{120'b111111111111111111111111111111101101111111111111111111101010111111111111111111111100000101111111111111111111111111110100},
{120'b011111111111111111111111111111101101111111111111111111010010111111111111111111111010000101111111111111111111111111101000},
{120'b011111111111111111111111111111101101111111111111111111010010111111111111111110101100000101111111111111111111111111100000},
{120'b101111111111111111111111111111101010111111111111111111010010111111111111111001111000000101111111111111111111111111010000},
{120'b101111111111111111111111111111010010111111111111111111010010111111111111101111111111111010111111111111111111111110100000},
{120'b010111111111111111111111111111010010111111111111111110100010111111111111111100000000000010111111111111111111111110100000},
{120'b010111111111111111111111111110100010111111111111111110100010111111111111111111111111111010111111111111111111111101000000},
{120'b001011111111111111111111111110100000011111111111111110100010111111111111111111111111111010111111111111111111111101000000},
{120'b001011111111111111111111111101000001011111111111111110100010111111111111111111111111111010111111111111111111111101000000},
{120'b000101111111111111111111111100000001011111111111111110100010111111111111111111111111111010111111111111111111111110100000},
{120'b000101111111111111111111111010000001011111111111111101000010111111111111111111111111111010111111111111111111111111011000},
{120'b000010111111111111111111110100000001011111111111111101000010111111111111111111111111111110111111111111111111111111101100},
{120'b000010111111111111111111110100000000101111111111111101000010111111111111111111111111111110111111111111111111111111111010},
{120'b000001011111111111111111101000000000101111111111111101000010111111111111111111111111111110111111111111111111111111111101},
{120'b000000001111111111111111101000000000101111111111111010000000011111111111111111111111111110111111111111111111111111111110},
{120'b000000101111111111111111010000000000101111111111111010000001011111111111111111111111111110111111111111111111111111111110},
{120'b000000010111111111111110100000000000010111111111111010000001011111111111111111111111111010111111111111111111111111111111},
{120'b000000000111111111111110100000000000010111111111111010000001011111111111111111111111111010111111111111111111111111111111},
{120'b000000000100000000000010000000000000010111111111111010000001011111111111111111111111111010111111111111111111111111111111},
{120'b000000000111111111111110000000000000010111111111110100000000011111111111111111111111111010111111111111011111111111111111},
{120'b000000000000000000000000000000000000001011111111110100000000000000000000000000000000000010111111111111001111111111111111},
{120'b000000000000000000000000000000000000001011111111110100000000001111111111111111111111111010111111111110110111111111111111},
{120'b000000000000000000000000000000000000001011111111110100000000000000000000000000000000000010111111111110101011111111111111},
{120'b000000000000000000000000000000000000001011111111101000000000000000000000000000000000000010111111111110100101111111111111},
{120'b000000000000000000000000000000000000000101111111101000000000000000000000000000000000000010111111111101000010111111111111},
{120'b000000000000000000000000000000000000000101111111101000000000000000000000000000000000000001011111111101000001000000000000}
};

int bCoord_X;// offset from start position 
int bCoord_Y;

logic drawing_X;
logic drawing_Y; // synthesis keep
logic mask_bit;
localparam int ObjectStartX = 260;
localparam int ObjectStartY = 180;
int objectEndX;
int objectEndY;



// Calculate object end boundaries
assign objectEndX    = (object_X_size + ObjectStartX);
assign objectEndY    = (object_Y_size + ObjectStartY);

// Signals drawing_X[Y] are active when obects coordinates are being crossed

// test if oCoord is in the rectangle defined by Start and End 
assign drawing_X  = ((oCoord_X  >= ObjectStartX) &&  (oCoord_X < objectEndX)) ? 1 : 0;
assign drawing_Y = ((oCoord_Y  >= ObjectStartY) &&  (oCoord_Y < objectEndY)) ? 1 : 0;

// calculate offset from start corner 
assign bCoord_X	= (drawing_X == 1 &&  drawing_Y == 1)  ? (oCoord_X - ObjectStartX): 0;
assign bCoord_Y	= (drawing_X == 1 &&  drawing_Y == 1  )  ? (oCoord_Y - ObjectStartY): 0; 


always_ff@ (posedge CLK, negedge RESETn)
begin
    if(!RESETn)
   begin
         mVGA_RGB	<= 8'b0;
         drawing_request     <= 1'b0;
         mask_bit	<=  1'b0;
    end
   else
  begin
			drawing_request	<= object_mask[bCoord_Y][bCoord_X] && drawing_X && drawing_Y && game_over_ena; // get from mask table if inside rectangle and enable
			mask_bit	<= object_mask[bCoord_Y][bCoord_X]; 
			if (object_mask[bCoord_Y][bCoord_X])
				mVGA_RGB <= 8'hE0; //uniform color
	end
end

endmodule		

//generated with PNGtoSV tool by Ben Wellingstein
